// Test
		// Test1

module example #( // here at the place
	parameter x = 5,
	// parameter
	parameter y = 4
)
(
	input clk,	// cent testing123
	output reg clk2,
	output reg [4:0] count,
	input [5 : 0] counter,
	input [ 6 : 0 ] counter_1,
	output reg [7: 0] counter_2

);

assign count = 1;


endmodule
