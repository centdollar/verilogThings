// Test
		// Test1

module example(
	input clk,
	output [4:0] count,
	input [4 : 0] counter,
	input [ 4 : 0 ] counter_1
);

assign count = 1;


endmodule
