// Test
		// Test1

module example #( // here at the place
	parameter x = 5,
	// parameter
	parameter y = 4
)
(
	input clk,	// cent Testing123
	output clk2,
	output [4:0] count,
	input [4 : 0] counter,
	input [ 4 : 0 ] counter_1,
	output [4: 0] counter_2

);

assign count = 1;


endmodule
